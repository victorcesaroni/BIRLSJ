LIBRARY ieee ;
	USE ieee.std_logic_1164.all;
	USE ieee.std_logic_signed.all;
	
ENTITY Projeto3 IS
	PORT(	CLOCK				: IN STD_LOGIC;
	
			DBG_PC 			: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_INSTRUCAO 	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			--DBG_PC_S1 		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			--DBG_INSTRUCAO_S1:OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			--DBG_OPCODE_S2	: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);			
			DBG_RegWrite_S4	: OUT STD_LOGIC;
			--DBG_ALUSrc		: OUT STD_LOGIC;
			--DBG_ALUOp		: OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
			--DBG_RegDst		: OUT STD_LOGIC;
			--DBG_MemWrite	: OUT STD_LOGIC;
			--DBG_MemRead		: OUT STD_LOGIC;
			--DBG_MemtoReg	: OUT STD_LOGIC;
			--DBG_PCSource 	: OUT STD_LOGIC;
			--DBG_Branch 		: OUT STD_LOGIC;
			--DBG_OPCODE 		: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			--DBG_FUNCT 		: OUT STD_LOGIC_VECTOR(5 DOWNTO 0)			
			
			DBG_REGWRITE_ADDR : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
			DBG_R0_DATA		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R1_DATA		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R2_DATA		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R3_DATA		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R4_DATA		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R5_DATA		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R6_DATA		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	) ;
END ENTITY ; -- Projeto3


ARCHITECTURE arch OF Projeto3 IS

	COMPONENT REGISTERS
		PORT(	CLOCK			: IN STD_LOGIC;
				REGWRITE		: IN STD_LOGIC;
				READ0_ADDR	: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
				READ1_ADDR	: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
				WRITE_ADDR 	: IN STD_LOGIC_VECTOR(4 DOWNTO 0);			
				WRITEDATA 	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				READ0_OUT 	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				READ1_OUT 	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			
				DBG_R0_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R1_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R2_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R3_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R4_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R5_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R6_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
	END COMPONENT; -- REGISTERS
	
	COMPONENT REG32
		GENERIC(N : INTEGER := 32);
		
		PORT(	CLOCK			: IN STD_LOGIC;
				ENTRADA 		: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
				REG_IN		: IN STD_LOGIC;
				SAIDA 		: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0) 
		);
	END COMPONENT; -- REG32
	
	COMPONENT REG32_DESCIDA
		GENERIC(N : INTEGER := 32);
		
		PORT(	CLOCK			: IN STD_LOGIC;
				ENTRADA 		: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
				REG_IN		: IN STD_LOGIC;
				SAIDA 		: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0) 
		);
	END COMPONENT; -- REG32_DESCIDA
	
	COMPONENT ADDER
		PORT(	ENTRADA_0 	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				ENTRADA_1	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				RESULT 		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
	END COMPONENT; -- ADDER
	
	COMPONENT MUX32_2_1
		PORT(	ENTRADA_0 	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				ENTRADA_1 	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				CONTROLE 	: IN STD_LOGIC;
				SAIDA 		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)		
		);
	END COMPONENT; -- MUX
	
	COMPONENT INSTRUCTIONMEMORY
		GENERIC(	N : INTEGER := 32 );
		
		PORT(	CLOCK 		: IN STD_LOGIC;
				PC				: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);				
				INSTRUCAO 	: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)
		);
	END COMPONENT; -- INSTRUCTIONMEMORY
	
	COMPONENT RegistradorIF_ID
		PORT( CLOCK		 	: IN STD_LOGIC;
				INSTRUCAO 	: IN STD_LOGIC_VECTOR(31 DOWNTO 0) ;
				PC			 	: IN STD_LOGIC_VECTOR(31 DOWNTO 0) ;				
				PC_OUT	 	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				INSTRUCAO_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
	END COMPONENT; -- RegistradorIF_ID
	
	COMPONENT DATAMEMORY IS
		GENERIC (N : INTEGER := 32);
				
		PORT(	CLOCK 		: IN STD_LOGIC;
				MEMWRITE 	: IN STD_LOGIC;
				MEMREAD		: IN STD_LOGIC;
				ADDRESS		: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
				WRITEDATA	: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
				READDATA		: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)
		);
	END COMPONENT; -- DATAMEMORY
	
	COMPONENT EXTENSOR IS  
		PORT( X 				: IN STD_LOGIC_VECTOR(18-1 DOWNTO 0) ;
				O 				: OUT STD_LOGIC_VECTOR(32-1 DOWNTO 0)
	);
	END COMPONENT; -- EXTENSOR
		
	COMPONENT RegistradorID_EX
	  PORT ( READ_DATA_1 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) ;
				READ_DATA_2 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) ;
				SINAL_EXTENDIDO : IN STD_LOGIC_VECTOR(31 DOWNTO 0) ; -- IMEDIATO
				RD			 	: IN STD_LOGIC_VECTOR(4 DOWNTO 0) ; -- RD
				PC			 	: IN STD_LOGIC_VECTOR(31 DOWNTO 0) ;
				OPCODE	 	: IN STD_LOGIC_VECTOR(3 DOWNTO 0) ;
				CLOCK		 	: IN STD_LOGIC;
				FUNCT 		: IN STD_LOGIC_VECTOR(5 DOWNTO 0);
				READ_DATA_1_OUT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				READ_DATA_2_OUT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				SINAL_EXTENDIDO_OUT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				RD_OUT		: OUT STD_LOGIC_VECTOR(4 DOWNTO 0) ; -- RD
				OPCODE_OUT	: OUT STD_LOGIC_VECTOR(3 DOWNTO 0); 
				PC_OUT	 	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				FUNCT_OUT	: OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
	  ) ;
	  
	END COMPONENT; -- RegistradorID_EX
	
	
	COMPONENT CONTROL
		PORT(	INSTRUCAO 	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				RegWrite		: OUT STD_LOGIC;
				ALUSrc		: OUT STD_LOGIC;
				ALUOp			: OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
				RegDst		: OUT STD_LOGIC;
				MemWrite		: OUT STD_LOGIC;
				MemRead		: OUT STD_LOGIC;
				MemtoReg		: OUT STD_LOGIC;
				Branch 		: OUT STD_LOGIC;
				OPCODE 		: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
				FUNCT 		: OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
		);
	END COMPONENT; -- CONTROL
	
	
	COMPONENT MUX32_3_1
		PORT(	ENTRADA_0 	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				ENTRADA_1 	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				ENTRADA_2 	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				CONTROLE 	: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
				SAIDA 		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)		
		);
	END COMPONENT; -- MUX
	
	COMPONENT RegistradorEX
	  PORT ( 	
				ALUSrc		: IN STD_LOGIC;
				ALUOp			: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
				RegDST		: IN STD_LOGIC;
				clock		 	: IN STD_LOGIC;
				ALUSrc_out	: OUT STD_LOGIC;
				ALUOp_out	: OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
				RegDST_out	: OUT STD_LOGIC				
	  );	  
	END COMPONENT; -- RegistradorEX
	
	
	COMPONENT RegistradorMEM
	  PORT ( 	
				MemWrite		: IN STD_LOGIC;
				MemRead		: IN STD_LOGIC;
				Branch		: IN STD_LOGIC;
				clock		 	: IN STD_LOGIC;
				MemWrite_out: OUT STD_LOGIC;
				MemRead_out	: OUT STD_LOGIC;
				Branch_out	: OUT STD_LOGIC
				
	  );	  
	END COMPONENT; -- RegistradorMEM
	
	COMPONENT RegistradorWB
	  PORT ( 	
				MemToReg		: IN STD_LOGIC;
				RegWrite		: IN STD_LOGIC;
				clock		 	: IN STD_LOGIC;
				MemToReg_out: OUT STD_LOGIC;
				RegWrite_out: OUT STD_LOGIC
				
	  );	  
	END COMPONENT; -- RegistradorWB
	
	COMPONENT RegistradorEX_MEM
	  PORT ( 	
				saidasomador			: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				sinalZero				: IN STD_LOGIC;
				ALUResult				: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				read_data_2 			: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				saida_mux_RegDST		: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
				clock		 				: IN STD_LOGIC;
				saidasomador_out		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				sinalZero_out			: OUT STD_LOGIC;
				ALUResult_out			: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				read_data_2_out		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				saida_mux_RegDST_out	: OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
	  );	  
	END COMPONENT; -- RegistradorEX_MEM	
	
	COMPONENT ALUControl  
	  PORT ( funct				: IN STD_LOGIC_VECTOR(5 DOWNTO 0) ;
				ALUOp 			: IN STD_LOGIC_VECTOR(2 DOWNTO 0) ;
				Opcode 			: IN STD_LOGIC_VECTOR(3 DOWNTO 0) ;
				operacao 		: OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
	  );
	END COMPONENT; -- ALUControl
	
	COMPONENT ALU
		PORT(	ALU_0 		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				ALU_1 		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				ALUOP 		: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
				RESULT 		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				ZERO 			: OUT STD_LOGIC
		);
	END COMPONENT; -- ALU
	
	COMPONENT MUX5_2_1
		PORT(	ENTRADA_0 	: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
				ENTRADA_1 	: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
				CONTROLE 	: IN STD_LOGIC;
				SAIDA 		: OUT STD_LOGIC_VECTOR(4 DOWNTO 0)		
		);
	END COMPONENT; -- MUX

	COMPONENT RegistradorMEM_WB
	  PORT ( 	
				read_data	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				address 		: IN STD_LOGIC_VECTOR(31 DOWNTO 0); -- CONFerir o tamanho
				saida_mux_RegDST: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
				clock		 	: IN STD_LOGIC;
				read_data_out:OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				address_out : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				saida_mux_RegDST_OUT: OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
	  );	  
	END COMPONENT; -- RegistradorMEM_WB

	SIGNAL READ0_ADDR		: STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL READ1_ADDR		: STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL RS_ADDR			: STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL RT_ADDR			: STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL RD_ADDR			: STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL REGWRITE_ADDR : STD_LOGIC_VECTOR(4 DOWNTO 0);			
	SIGNAL REGWRITEDATA 	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL REG0_DATA 		: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL REG1_DATA 		: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL PC_DATA 		: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL PC_MAIS_UM		: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL PC_PROX			: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL PC_BRANCH 		: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL PC_REG	 		: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL INSTRUCAO 		: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL INSTRUCAO_S1	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL PC_S1 			: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL IMMED_EXT 		: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL REG0_DATA_S2	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL REG1_DATA_S2	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL IMMED_EXT_S2	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL RD_ADDR_S2		: STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL OPCODE_S2		: STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL PC_S2 			: STD_LOGIC_VECTOR(31 DOWNTO 0);

	SIGNAL MEMADDRESS 	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL MEMWRITE_DATA	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL MEMREAD_DATA 	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	
	SIGNAL RegWrite		: STD_LOGIC;
	SIGNAL ALUSrc			: STD_LOGIC;
	SIGNAL ALUOp			: STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL RegDst			: STD_LOGIC;
	SIGNAL MemWrite		: STD_LOGIC;
	SIGNAL MemRead			: STD_LOGIC;
	SIGNAL MemtoReg		: STD_LOGIC;
	SIGNAL PCSource_S3 	: STD_LOGIC;	
	SIGNAL Branch 			: STD_LOGIC;
	SIGNAL OPCODE 			: STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL FUNCT 			: STD_LOGIC_VECTOR(5 DOWNTO 0);	
	
	SIGNAL ALUSrc_S2		: STD_LOGIC;
	SIGNAL ALUOp_S2		: STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL RegDst_S2		: STD_LOGIC;
	
	SIGNAL MemWrite_S2 	: STD_LOGIC;
	SIGNAL MemRead_S2		: STD_LOGIC;
	SIGNAL Branch_S2		: STD_LOGIC;
	
	SIGNAL MemToReg_S2	: STD_LOGIC;
	SIGNAL RegWrite_S2	: STD_LOGIC;
	
	SIGNAL MemWrite_S3 	: STD_LOGIC;
	SIGNAL MemRead_S3		: STD_LOGIC;
	SIGNAL Branch_S3		: STD_LOGIC;
	
	SIGNAL MemToReg_S3	: STD_LOGIC;
	SIGNAL RegWrite_S3	: STD_LOGIC;
	
	SIGNAL MemToReg_S4	: STD_LOGIC;
	SIGNAL RegWrite_S4	: STD_LOGIC;	
	
	SIGNAL SOMADOR			: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL ZERO				: STD_LOGIC;
	SIGNAL ALUResult		: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL REG1_DATA_S3 	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL REGDST_S3		: STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL SOMADOR_S3		: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL ZERO_S3			: STD_LOGIC;
	SIGNAL ALUResult_S3	: STD_LOGIC_VECTOR(31 DOWNTO 0);

	SIGNAL FUNCT_S2 		: STD_LOGIC_VECTOR(5 DOWNTO 0);

	SIGNAL OPERACAO_ALU_S2:STD_LOGIC_VECTOR(2 DOWNTO 0);
	
	SIGNAL ALU_0_S2 		: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL ALU_1_S2 		: STD_LOGIC_VECTOR(31 DOWNTO 0);
	
	SIGNAL MUX_REG_DST_S2: STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL MUX_REG_DST_S3: STD_LOGIC_VECTOR(4 DOWNTO 0);
	
	SIGNAL MEMREAD_DATA_S3:STD_LOGIC_VECTOR(31 DOWNTO 0);
	
	SIGNAL MEMREAD_DATA_S4:STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL ADDRESS_S4		: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL MUX_REG_DST_S4: STD_LOGIC_VECTOR(4 DOWNTO 0);
	
	SIGNAL RegWriteAddr_S4:STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL RegWriteData_S4:STD_LOGIC_VECTOR(31 DOWNTO 0);
	

BEGIN
	
	-- TESTE TESTE TESTE TESTE TESTE
	--PCSOURCE <= '0';
	--PC_BRANCH <= "01010101010101010101010101010101";
	--------------------------------

	-------------------------------------------------------------------------------------------
	-- IF 1
	PC0: REG32_DESCIDA PORT MAP(	
				CLOCK, 
				PC_PROX, 
				'1', 
				PC_DATA
	);
								
	ADDERPC0: ADDER PORT MAP(	
				PC_DATA, 
				"00000000000000000000000000000001",	
				PC_MAIS_UM
	);
										
	MUXPC0: MUX32_2_1 PORT MAP(
				PC_MAIS_UM, 
				PC_BRANCH, 
				PCSOURCE_S3,
				PC_PROX
	);	
	
	INSTRUCTIONMEMORY0: INSTRUCTIONMEMORY PORT MAP(	
				CLOCK, 
				PC_DATA, 
				INSTRUCAO
	);
	
	RegistradorIF_ID0: RegistradorIF_ID PORT MAP(	
				CLOCK, 
				INSTRUCAO, 
				PC_MAIS_UM,
				PC_S1, 
				INSTRUCAO_S1
	);
																
	-------------------------------------------------------------------------------------------
	-- ID 2
	RD_ADDR <= INSTRUCAO_S1(27 DOWNTO 23); -- rd
	RS_ADDR <= INSTRUCAO_S1(22 DOWNTO 18); -- rs	
	RT_ADDR <= INSTRUCAO_S1(17 DOWNTO 13); -- rt
	
	REGWRITE_ADDR <= RegWriteAddr_S4;
	
	EXTENSORIMMED0: EXTENSOR PORT MAP(
				INSTRUCAO_S1(17 DOWNTO 0), 
				IMMED_EXT
	);	
	
	REGISTERS0: REGISTERS PORT MAP(	
				CLOCK, 
				RegWrite_S4, 
				RS_ADDR, 
				RT_ADDR, 
				REGWRITE_ADDR, 
				RegWriteData_S4,
				REG0_DATA, 
				REG1_DATA,
				DBG_R0_DATA,
				DBG_R1_DATA,
				DBG_R2_DATA,
				DBG_R3_DATA,
				DBG_R4_DATA,
				DBG_R5_DATA,
				DBG_R6_DATA
	);
											
	CONTROL0: CONTROL PORT MAP(	INSTRUCAO_S1, 
				RegWrite, 
				ALUSrc,
				ALUOp,
				RegDst,
				MemWrite,
				MemRead,
				MemtoReg,
				Branch,
				OPCODE, 
				FUNCT 
	);
	
	RegistradorID_EX0: RegistradorID_EX PORT MAP(
				REG0_DATA, 
				REG1_DATA, 
				IMMED_EXT,
				RD_ADDR,
				PC_S1,
				OPCODE,
				CLOCK,
				INSTRUCAO_S1(5 DOWNTO 0),
				REG0_DATA_S2,
				REG1_DATA_S2,
				IMMED_EXT_S2,
				RD_ADDR_S2,
				OPCODE_S2,
				PC_S2,
				FUNCT_S2);
			
			
	RegistradorEX_0: RegistradorEX PORT MAP(
				ALUSrc,
				ALUOp,		
				RegDst,
				CLOCK,
				ALUSrc_S2,	
				ALUOp_S2,	
				RegDST_S2			
	);
	
	
	RegistradorMEM_0: RegistradorMEM PORT MAP(
				MemWrite,
				MemRead,
				Branch,
				CLOCK,
				MemWrite_S2,
				MemRead_S2,
				Branch_S2
	);
	
	RegistradorWB_0: RegistradorWB PORT MAP(	  
				MemToReg,
				RegWrite,
				CLOCK,
				MemToReg_S2,
				RegWrite_S2		
	);
	
	-------------------------------------------------------------------------------------------
	-- EX 3
		
	MUXALU0: MUX32_2_1 PORT MAP(
				REG1_DATA_S2,
				IMMED_EXT_S2,
				ALUSrc_S2,
				ALU_1_S2				
	);	
	
	-- MUX nao necessario, alterar depois
	MUXREGDST: MUX5_2_1 PORT MAP(
				RD_ADDR_S2,
				RD_ADDR_S2,
				REGDST_S2,
				MUX_REG_DST_S2
	);	


	RegistradorEX_MEM0: RegistradorEX_MEM PORT MAP(
				SOMADOR,
				ZERO,
				ALUResult,
				REG1_DATA_S2,
				MUX_REG_DST_S2,
				CLOCK,
				SOMADOR_S3,
				ZERO_S3,
				ALUResult_S3,
				REG1_DATA_S3,
				MUX_REG_DST_S3
	);
	
	
	ALUControl0: ALUControl PORT MAP(
				FUNCT_S2,
				ALUOp_S2,
				OPCODE_S2,
				OPERACAO_ALU_S2
	);
	
	ALU0: ALU PORT MAP(
				ALU_0_S2,
				ALU_1_S2,
				OPERACAO_ALU_S2,
				ALUResult,
				ZERO
	);
	
	ADDERBRANCH0: ADDER PORT MAP(	
				PC_S2, 
				IMMED_EXT_S2,	
				SOMADOR
	);
	
	RegistradorMEM_1: RegistradorMEM PORT MAP(
				MemWrite_S2,
				MemRead_S2,
				Branch_S2,
				CLOCK,
				MemWrite_S3,
				MemRead_S3,
				Branch_S3
	);
	
	RegistradorWB_1: RegistradorWB PORT MAP(	  
				MemToReg_S2,
				RegWrite_S2,
				CLOCK,
				MemToReg_S3,
				RegWrite_S3		
	);
	
		
	-------------------------------------------------------------------------------------------
	-- MEM 4
	DATAMEMORY0: DATAMEMORY PORT MAP(	
				CLOCK, 
				MEMWRITE_S3, 
				MEMREAD_S3,
				ALUResult_S3, 
				REG1_DATA_S3, 
				MEMREAD_DATA_S3
	);	
	
	PCSource_S3 <= Branch AND ZERO_S3;
	
	RegistradorMEM_WB0: RegistradorMEM_WB PORT MAP(
				MEMREAD_DATA_S3,
				ALUResult_S3,
				MUX_REG_DST_S3,
				CLOCK,
				MEMREAD_DATA_S4,
				ADDRESS_S4,
				MUX_REG_DST_S4
	);
	
	RegistradorWB_2: RegistradorWB PORT MAP(	  
				MemToReg_S3,
				RegWrite_S3,
				CLOCK,
				MemToReg_S4,
				RegWrite_S4		
	);

	
	-------------------------------------------------------------------------------------------
	-- WB	5
	
	RegWriteAddr_S4 <= MUX_REG_DST_S4;
		
	MUXMEMTOREG: MUX32_2_1 PORT MAP(
				ADDRESS_S4,
				IMMED_EXT_S2,
				MemToReg_S4,
				RegWriteData_S4	
	);	
	

	-------------------------------------------------------------------------------------------
	-- DBG
	
	DBG_REGWRITE_ADDR <= REGWRITE_ADDR;
	DBG_PC <= PC_DATA;
	DBG_INSTRUCAO <= INSTRUCAO;
	--DBG_PC_S1 <= PC_S1;
	--DBG_INSTRUCAO_S1 <= INSTRUCAO_S1;
	--DBG_OPCODE_S2 <= OPCODE_S2;
	
	DBG_RegWrite_S4	<= RegWrite_S4;
	--DBG_ALUSrc		<= ALUSrc;
	--DBG_ALUOp		<= ALUOp;
	--DBG_RegDst		<= RegDst;
	--DBG_MemWrite	<= MemWrite;
	--DBG_MemRead		<= MemRead;
	--DBG_MemtoReg	<= MemtoReg;
	--DBG_PCSource 	<= PCSource_S3;
	--DBG_Branch 		<= Branch;
	--DBG_OPCODE 		<= OPCODE; 	
	--DBG_FUNCT 		<= FUNCT;
	
END ARCHITECTURE ; -- arch