LIBRARY ieee ;
USE ieee.std_logic_1164.all ;

ENTITY REG32 IS
	GENERIC(N : INTEGER := 32);
	
	PORT(	CLOCK		: IN STD_LOGIC;
			ENTRADA 	: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
			REG_IN	: IN STD_LOGIC;
			SAIDA 	: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0) 
	);
END REG32 ;


ARCHITECTURE Behavior OF REG32 IS
BEGIN
	PROCESS (CLOCK, REG_IN)
	BEGIN
		IF (CLOCK'EVENT AND CLOCK = '1') THEN		
			IF REG_IN = '1' THEN
				SAIDA <= ENTRADA;
			END IF ;
		END IF;
	END PROCESS ;
END Behavior ;
