library ieee ;
	use ieee.std_logic_1164.all ;
	use ieee.numeric_std.all ;

ENTITY MUX32_3_1 IS
	PORT(	ENTRADA_0 	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			ENTRADA_1 	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			ENTRADA_2 	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			CONTROLE 	: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
			SAIDA 		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)		
	) ;
END ENTITY ; -- MUX

ARCHITECTURE arch OF MUX32_3_1 IS
BEGIN
	PROCESS (CONTROLE, ENTRADA_0, ENTRADA_1, ENTRADA_2)
		BEGIN
		CASE CONTROLE IS
			WHEN "00" => SAIDA <= ENTRADA_0;
			WHEN "01" => SAIDA <= ENTRADA_1;
			WHEN "10" => SAIDA <= ENTRADA_2;
			WHEN OTHERS => NULL;
		END CASE;
	END PROCESS;
END ARCHITECTURE ; -- arch