LIBRARY ieee ;
	USE ieee.std_logic_1164.all;
	USE ieee.std_logic_signed.all;
	USE ieee.numeric_std.all;
	
ENTITY REGISTERS IS
	GENERIC(	N : INTEGER := 32; 
				M : INTEGER := 32
	); -- registradores de 32bits x 32
	
	
	PORT(	CLOCK			: IN STD_LOGIC;
			REGWRITE		: IN STD_LOGIC;
			READ0_ADDR	: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			READ1_ADDR	: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			WRITE_ADDR 	: IN STD_LOGIC_VECTOR(4 DOWNTO 0);			
			WRITEDATA 	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			READ0_OUT 	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			READ1_OUT 	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	
			DBG_R0_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R1_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R2_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R3_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R4_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R5_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R6_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R7_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R8_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R9_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R10_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R11_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R12_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R13_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R14_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R15_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R16_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R17_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R18_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R19_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R20_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R21_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R22_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R23_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R24_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R25_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R26_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R27_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R28_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R29_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R30_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R31_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	) ;
END ENTITY ; -- REGISTERS


ARCHITECTURE arch OF REGISTERS IS
	TYPE REGISTERS_ARRAY IS ARRAY (0 TO M-1) OF STD_LOGIC_VECTOR(N-1 DOWNTO 0);	
	SIGNAL REGS : REGISTERS_ARRAY;	
	
	SIGNAL READ0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL READ1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
		
BEGIN
	
	PROCESS (CLOCK)
	BEGIN
		IF (CLOCK'EVENT AND CLOCK = '1') THEN
			IF(REGWRITE = '1') THEN
				REGS(TO_INTEGER(UNSIGNED(WRITE_ADDR))) <= WRITEDATA;
			END IF;
		END IF;
		
		READ0 <= REGS(TO_INTEGER(UNSIGNED(READ0_ADDR)));
		READ1 <= REGS(TO_INTEGER(UNSIGNED(READ1_ADDR)));
	END PROCESS;
		
	READ0_OUT <= READ0;
	READ1_OUT <= READ1;
	
	DBG_R0_DATA <= REGS(0);
	DBG_R1_DATA <= REGS(1);
	DBG_R2_DATA <= REGS(2);
	DBG_R3_DATA <= REGS(3);
	DBG_R4_DATA <= REGS(4);
	DBG_R5_DATA <= REGS(5);
	DBG_R6_DATA <= REGS(6);
	DBG_R7_DATA <= REGS(7);
	DBG_R8_DATA <= REGS(8);
	DBG_R9_DATA <= REGS(9);
	DBG_R10_DATA<= REGS(10);
	DBG_R11_DATA<= REGS(11);
	DBG_R12_DATA<= REGS(12);
	DBG_R13_DATA<= REGS(13);
	DBG_R14_DATA<= REGS(14);
	DBG_R15_DATA<= REGS(15);
	DBG_R16_DATA<= REGS(16);
	DBG_R17_DATA<= REGS(17);
	DBG_R18_DATA<= REGS(18);
	DBG_R19_DATA<= REGS(19);
	DBG_R20_DATA<= REGS(20);
	DBG_R21_DATA<= REGS(21);
	DBG_R22_DATA<= REGS(22);
	DBG_R23_DATA<= REGS(23);
	DBG_R24_DATA<= REGS(24);
	DBG_R25_DATA<= REGS(25);
	DBG_R26_DATA<= REGS(26);
	DBG_R27_DATA<= REGS(27);
	DBG_R28_DATA<= REGS(28);
	DBG_R29_DATA<= REGS(29);
	DBG_R30_DATA<= REGS(30);
	DBG_R31_DATA<= REGS(31);
	
END ARCHITECTURE ; -- arch