LIBRARY ieee ;
	USE ieee.std_logic_1164.all;
	USE ieee.std_logic_signed.all;
	
ENTITY Projeto3_V2 IS
	PORT(	CLOCK					: IN STD_LOGIC;
	
			DBG_PC_IF			: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			--DBG_PC_ID			: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_INSTRUCAO_IF 	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			--DBG_INSTRUCAO_ID	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);			
						
			--DBG_REGWRITE_ID	: OUT STD_LOGIC;
			--DBG_REGWRITE_EX	: OUT STD_LOGIC;
			--DBG_REGWRITE_MEM 	: OUT STD_LOGIC;
			
			--DBG_RegWrite_WB 		: OUT STD_LOGIC;
			--DBG_RD_ADDR_WB 		: OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
			--DBG_RegWriteData_WB 	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			--DBG_MEMREAD_DATA_WB	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			--DBG_ALUResult_WB		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			--DBG_MemToReg_WB		: OUT  STD_LOGIC;
			
			--DBG_RS_DATA_ID		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			--DBG_RT_DATA_ID		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			--DBG_RS_ADDR_ID 	: OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
			--DBG_RT_ADDR_ID 	: OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
			
			--DBG_RS_DATA_EX		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			--DBG_RT_DATA_EX		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			
			--DBG_OPERACAO_ALU_EX 	: OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
			--DBG_FUNCT_EX 		: OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
			
			--DBG_MemWrite_MEM 	: OUT STD_LOGIC;
			--DBG_MemRead_MEM 	: OUT STD_LOGIC;
			--DBG_ALUResult_MEM : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			--DBG_RT_DATA_MEM 	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			
			--DBG_Branch_MEM 	: OUT STD_LOGIC;
			--DBG_ZERO_MEM 		: OUT STD_LOGIC;
			--DBG_SOMADOR_MEM 	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			
			DBG_R0_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R1_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R2_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R3_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R4_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R5_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R6_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R7_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R8_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R9_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R10_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R11_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R12_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R13_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R14_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R15_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R16_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R17_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R18_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R19_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R20_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R21_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R22_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R23_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R24_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R25_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R26_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R27_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R28_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R29_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R30_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DBG_R31_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);

			
			DBG_MEM0		: out std_logic_vector(31 downto 0);
			DBG_MEM1		: out std_logic_vector(31 downto 0);
			DBG_MEM2		: out std_logic_vector(31 downto 0);
			DBG_MEM3		: out std_logic_vector(31 downto 0);
			DBG_MEM4		: out std_logic_vector(31 downto 0);
			DBG_MEM5		: out std_logic_vector(31 downto 0);
			DBG_MEM6		: out std_logic_vector(31 downto 0);
			DBG_MEM7		: out std_logic_vector(31 downto 0)
	) ;
END ENTITY ; -- Projeto3_V2


ARCHITECTURE arch OF Projeto3_V2 IS

	COMPONENT REGISTERS
		PORT(	CLOCK			: IN STD_LOGIC;
				REGWRITE		: IN STD_LOGIC;
				READ0_ADDR	: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
				READ1_ADDR	: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
				WRITE_ADDR 	: IN STD_LOGIC_VECTOR(4 DOWNTO 0);			
				WRITEDATA 	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				READ0_OUT 	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				READ1_OUT 	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			
				DBG_R0_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R1_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R2_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R3_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R4_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R5_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R6_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R7_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R8_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R9_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R10_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R11_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R12_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R13_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R14_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R15_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R16_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R17_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R18_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R19_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R20_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R21_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R22_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R23_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R24_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R25_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R26_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R27_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R28_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R29_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R30_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				DBG_R31_DATA: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
	END COMPONENT; -- REGISTERS
	
	COMPONENT REG32
		GENERIC(N : INTEGER := 32);
		
		PORT(	CLOCK			: IN STD_LOGIC;
				ENTRADA 		: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
				REG_IN		: IN STD_LOGIC;
				SAIDA 		: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0) 
		);
	END COMPONENT; -- REG32
	
	COMPONENT REG32_DESCIDA
		GENERIC(N : INTEGER := 32);
		
		PORT(	CLOCK			: IN STD_LOGIC;
				ENTRADA 		: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
				REG_IN		: IN STD_LOGIC;
				SAIDA 		: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0) 
		);
	END COMPONENT; -- REG32_DESCIDA
	
	COMPONENT ADDER
		PORT(	ENTRADA_0 	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				ENTRADA_1	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				RESULT 		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
	END COMPONENT; -- ADDER
	
	COMPONENT MUX32_2_1
		PORT(	ENTRADA_0 	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				ENTRADA_1 	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				CONTROLE 	: IN STD_LOGIC;
				SAIDA 		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)		
		);
	END COMPONENT; -- MUX
	
	COMPONENT INSTRUCTIONMEMORY
		GENERIC(	N : INTEGER := 32 );
		
		PORT(	CLOCK 		: IN STD_LOGIC;
				PC				: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);				
				INSTRUCAO 	: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)
		);
	END COMPONENT; -- INSTRUCTIONMEMORY
	
	COMPONENT RegistradorIF_ID
		PORT( CLOCK		 	: IN STD_LOGIC;
				INSTRUCAO 	: IN STD_LOGIC_VECTOR(31 DOWNTO 0) ;
				PC			 	: IN STD_LOGIC_VECTOR(31 DOWNTO 0) ;				
				PC_OUT	 	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				INSTRUCAO_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
	END COMPONENT; -- RegistradorIF_ID
	
	COMPONENT DATAMEMORY IS
		GENERIC (N : INTEGER := 32);
				
		PORT(	CLOCK 		: IN STD_LOGIC;
				MEMWRITE 	: IN STD_LOGIC;
				MEMREAD		: IN STD_LOGIC;
				ADDRESS		: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
				WRITEDATA	: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
				READDATA		: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0);
				
				DBG_MEM0		: out std_logic_vector(N-1 downto 0);
				DBG_MEM1		: out std_logic_vector(N-1 downto 0);
				DBG_MEM2		: out std_logic_vector(N-1 downto 0);
				DBG_MEM3		: out std_logic_vector(N-1 downto 0);
				DBG_MEM4		: out std_logic_vector(N-1 downto 0);
				DBG_MEM5		: out std_logic_vector(N-1 downto 0);
				DBG_MEM6		: out std_logic_vector(N-1 downto 0);
				DBG_MEM7		: out std_logic_vector(N-1 downto 0)
		);
	END COMPONENT; -- DATAMEMORY
	
	COMPONENT EXTENSOR IS  
		PORT( X 				: IN STD_LOGIC_VECTOR(18-1 DOWNTO 0) ;
				O 				: OUT STD_LOGIC_VECTOR(32-1 DOWNTO 0)
	);
	END COMPONENT; -- EXTENSOR
		
	COMPONENT RegistradorID_EX
	  PORT ( READ_DATA_1 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) ;
				READ_DATA_2 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) ;
				SINAL_EXTENDIDO : IN STD_LOGIC_VECTOR(31 DOWNTO 0) ; -- IMEDIATO
				RD			 	: IN STD_LOGIC_VECTOR(4 DOWNTO 0) ; -- RD
				PC			 	: IN STD_LOGIC_VECTOR(31 DOWNTO 0) ;
				OPCODE	 	: IN STD_LOGIC_VECTOR(3 DOWNTO 0) ;
				CLOCK		 	: IN STD_LOGIC;
				FUNCT 		: IN STD_LOGIC_VECTOR(5 DOWNTO 0);
				READ_DATA_1_OUT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				READ_DATA_2_OUT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				SINAL_EXTENDIDO_OUT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				RD_OUT		: OUT STD_LOGIC_VECTOR(4 DOWNTO 0) ; -- RD
				OPCODE_OUT	: OUT STD_LOGIC_VECTOR(3 DOWNTO 0); 
				PC_OUT	 	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				FUNCT_OUT	: OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
	  ) ;
	  
	END COMPONENT; -- RegistradorID_EX
	
	
	COMPONENT CONTROL
		PORT(
				CLOCK			: IN STD_LOGIC;
				INSTRUCAO 	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				RegWrite		: OUT STD_LOGIC;
				ALUSrc		: OUT STD_LOGIC;
				ALUOp			: OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
				RegDst		: OUT STD_LOGIC;
				MemWrite		: OUT STD_LOGIC;
				MemRead		: OUT STD_LOGIC;
				MemtoReg		: OUT STD_LOGIC;
				Branch 		: OUT STD_LOGIC;
				OPCODE 		: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
				FUNCT 		: OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
				RD_ADDR		: OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
				RS_ADDR		: OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
				RT_ADDR		: OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
				AddSrc 		: OUT STD_LOGIC;
				Jump			: OUT STD_LOGIC;
				ImmedOrReg 	: OUT STD_LOGIC
		);
	END COMPONENT; -- CONTROL
	
	
	COMPONENT MUX32_3_1
		PORT(	ENTRADA_0 	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				ENTRADA_1 	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				ENTRADA_2 	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				CONTROLE 	: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
				SAIDA 		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)		
		);
	END COMPONENT; -- MUX
	
	COMPONENT RegistradorEX
	  PORT ( 	
				ALUSrc		: IN STD_LOGIC;
				ALUOp			: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
				RegDST		: IN STD_LOGIC;
				clock		 	: IN STD_LOGIC;
				AddSrc 		: IN STD_LOGIC;	
				ImmedOrReg	: IN STD_LOGIC;
				ALUSrc_out	: OUT STD_LOGIC;
				ALUOp_out	: OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
				RegDST_out	: OUT STD_LOGIC;
				AddSrc_out 	: OUT STD_LOGIC;
				ImmedOrReg_out:OUT STD_LOGIC
	  );	  
	END COMPONENT; -- RegistradorEX
	
	
	COMPONENT RegistradorMEM
	  PORT ( 	
				MemWrite		: IN STD_LOGIC;
				MemRead		: IN STD_LOGIC;
				Branch		: IN STD_LOGIC;
				clock		 	: IN STD_LOGIC;
				Jump 			: IN STD_LOGIC;
				MemWrite_out: OUT STD_LOGIC;
				MemRead_out	: OUT STD_LOGIC;
				Branch_out	: OUT STD_LOGIC;
				Jump_out 	: OUT STD_LOGIC
				
	  );	  
	END COMPONENT; -- RegistradorMEM
	
	COMPONENT RegistradorWB
	  PORT ( 	
				MemToReg		: IN STD_LOGIC;
				RegWrite		: IN STD_LOGIC;
				clock		 	: IN STD_LOGIC;
				MemToReg_out: OUT STD_LOGIC;
				RegWrite_out: OUT STD_LOGIC
				
	  );	  
	END COMPONENT; -- RegistradorWB
	
	COMPONENT RegistradorEX_MEM
	  PORT ( 	
				saidasomador			: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				sinalZero				: IN STD_LOGIC;
				ALUResult				: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				read_data_2 			: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				saida_mux_RegDST		: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
				clock		 				: IN STD_LOGIC;
				saidasomador_out		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				sinalZero_out			: OUT STD_LOGIC;
				ALUResult_out			: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				read_data_2_out		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				saida_mux_RegDST_out	: OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
	  );	  
	END COMPONENT; -- RegistradorEX_MEM	
	
	COMPONENT ALUControl  
	  PORT ( funct				: IN STD_LOGIC_VECTOR(5 DOWNTO 0) ;
				ALUOp 			: IN STD_LOGIC_VECTOR(2 DOWNTO 0) ;
				Opcode 			: IN STD_LOGIC_VECTOR(3 DOWNTO 0) ;
				operacao 		: OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
	  );
	END COMPONENT; -- ALUControl
	
	COMPONENT ALU
		PORT(	ALU_0 		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				ALU_1 		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				ALUOP 		: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
				RESULT 		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				ZERO 			: OUT STD_LOGIC
		);
	END COMPONENT; -- ALU
	
	COMPONENT MUX5_2_1
		PORT(	ENTRADA_0 	: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
				ENTRADA_1 	: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
				CONTROLE 	: IN STD_LOGIC;
				SAIDA 		: OUT STD_LOGIC_VECTOR(4 DOWNTO 0)		
		);
	END COMPONENT; -- MUX

	COMPONENT RegistradorMEM_WB
	  PORT ( 	
				read_data	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				address 		: IN STD_LOGIC_VECTOR(31 DOWNTO 0); -- CONFerir o tamanho
				saida_mux_RegDST: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
				clock		 	: IN STD_LOGIC;
				read_data_out:OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				address_out : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				saida_mux_RegDST_OUT: OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
	  );	  
	END COMPONENT; -- RegistradorMEM_WB
	
	SIGNAL PC_IF			: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL PC_PROX_IF		: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL PC_MAIS_UM_IF	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL INSTRUCAO_IF 	: STD_LOGIC_VECTOR(31 DOWNTO 0);	
	
	SIGNAL PC_ID 			: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL INSTRUCAO_ID 	: STD_LOGIC_VECTOR(31 DOWNTO 0);	
	SIGNAL FUNCT_ID 		: STD_LOGIC_VECTOR(5 DOWNTO 0);
	SIGNAL RegWrite_ID	: STD_LOGIC;
	SIGNAL ALUSrc_ID		: STD_LOGIC;	
	SIGNAL ALUOp_ID		: STD_LOGIC_VECTOR(2 DOWNTO 0);	
	SIGNAL RegDst_ID		: STD_LOGIC;
	SIGNAL MemWrite_ID	: STD_LOGIC;
	SIGNAL MemRead_ID		: STD_LOGIC;
	SIGNAL MemtoReg_ID	: STD_LOGIC;
	SIGNAL Branch_ID		: STD_LOGIC;
	SIGNAL OPCODE_ID		: STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL RD_ADDR_ID 	: STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL RS_ADDR_ID 	: STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL RT_ADDR_ID 	: STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL AddSrc_ID 		: STD_LOGIC;
	SIGNAL Jump_ID 		: STD_LOGIC;
	SIGNAL ImmedOrReg_ID	: STD_LOGIC;

	SIGNAL PCSource_MEM 	: STD_LOGIC;
	
	SIGNAL IMMED_EXT_ID 	: STD_LOGIC_VECTOR(31 DOWNTO 0);	
	SIGNAL RS_DATA_ID 	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL RT_DATA_ID 	: STD_LOGIC_VECTOR(31 DOWNTO 0);

	SIGNAL RS_DATA_EX		: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL RT_DATA_EX		: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL IMMED_EXT_EX	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL RD_ADDR_EX 	: STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL OPCODE_EX		: STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL PC_EX			: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL FUNCT_EX		: STD_LOGIC_VECTOR(5 DOWNTO 0);
	SIGNAL ALUSrc_EX	 	: STD_LOGIC;
	SIGNAL ALUOp_EX		: STD_LOGIC_VECTOR(2 DOWNTO 0);	
	SIGNAL RegDST_EX		: STD_LOGIC;
	SIGNAL MemWrite_EX	: STD_LOGIC;
	SIGNAL MemRead_EX 	: STD_LOGIC;
	SIGNAL Branch_EX		: STD_LOGIC;
	SIGNAL MemToReg_EX 	: STD_LOGIC;
	SIGNAL RegWrite_EX 	: STD_LOGIC;
	SIGNAL ALU_B_EX		: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL SOMADOR_EX		: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL OPERACAO_ALU_EX:STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL ALUResult_EX	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL ZERO_EX			: STD_LOGIC;
	SIGNAL AddSrc_EX 		: STD_LOGIC;
	SIGNAL Jump_EX 		: STD_LOGIC;
	SIGNAL ADDER_A_EX 	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL ImmedOrReg_EX	: STD_LOGIC;
	SIGNAL SOMADOR_TMP_EX: STD_LOGIC_VECTOR(31 DOWNTO 0);
	
	SIGNAL SOMADOR_MEM	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL ZERO_MEM		: STD_LOGIC;
	SIGNAL ALUResult_MEM	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL RT_DATA_MEM	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL RD_ADDR_MEM	: STD_LOGIC_VECTOR(4 DOWNTO 0);	
	SIGNAL MemWrite_MEM 	: STD_LOGIC;
	SIGNAL MemRead_MEM	: STD_LOGIC;
	SIGNAL Branch_MEM		: STD_LOGIC;
	SIGNAL MemToReg_MEM	: STD_LOGIC;
	SIGNAL RegWrite_MEM	: STD_LOGIC;
	SIGNAL MEMREAD_DATA_MEM	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL Jump_MEM 		: STD_LOGIC;	
			
	SIGNAL RegWrite_WB 		: STD_LOGIC;
	SIGNAL RD_ADDR_WB 		: STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL RegWriteData_WB 	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL MEMREAD_DATA_WB	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL ALUResult_WB		: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL MemToReg_WB		: STD_LOGIC;


BEGIN
	

	-------------------------------------------------------------------------------------------
	-- IF 1
	
	-- REG PC
	PC0: REG32_DESCIDA PORT MAP(
				-- in
				CLOCK, 
				PC_PROX_IF, 
				'1',
				-- out
				PC_IF
	);
	
	-- PC + 1
	ADDERPC0: ADDER PORT MAP(	
				-- in
				PC_IF, 
				"00000000000000000000000000000001",	
				-- out
				PC_MAIS_UM_IF
	);
	
	-- PCSource MUX
	MUXPC0: MUX32_2_1 PORT MAP(
				-- in
				PC_MAIS_UM_IF, 
				SOMADOR_MEM, 
				PCSource_MEM,
				-- out
				PC_PROX_IF
	);
	
	-- INSTRUCTION MEMORY
	INSTRUCTIONMEMORY0: INSTRUCTIONMEMORY PORT MAP(	
				--in
				CLOCK, 
				PC_IF,				
				-- out
				INSTRUCAO_IF
	);
	
	-- REG PIPELINE IF/ID	
	RegistradorIF_ID0: RegistradorIF_ID PORT MAP(	
				-- in
				CLOCK, 
				INSTRUCAO_IF, 
				PC_IF,
				-- out
				PC_ID, 
				INSTRUCAO_ID
	);
																
	-------------------------------------------------------------------------------------------
	-- ID 2
	
	-- Extensor de sinal
	EXTENSORIMMED0: EXTENSOR PORT MAP(
				-- in
				INSTRUCAO_ID(17 DOWNTO 0), 
				-- out
				IMMED_EXT_ID
	);	
	
	
	-- Banco de Registradores
	REGISTERS0: REGISTERS PORT MAP(
				-- in
				CLOCK, 
				RegWrite_WB, 
				RS_ADDR_ID, 
				RT_ADDR_ID, 
				RD_ADDR_WB, 
				RegWriteData_WB,
				-- out
				RS_DATA_ID, 
				RT_DATA_ID,
				DBG_R0_DATA,
				DBG_R1_DATA,
				DBG_R2_DATA,
				DBG_R3_DATA,
				DBG_R4_DATA,
				DBG_R5_DATA,
				DBG_R6_DATA,
				DBG_R7_DATA,
				DBG_R8_DATA,
				DBG_R9_DATA,
				DBG_R10_DATA,
				DBG_R11_DATA,
				DBG_R12_DATA,
				DBG_R13_DATA,
				DBG_R14_DATA,
				DBG_R15_DATA,
				DBG_R16_DATA,
				DBG_R17_DATA,
				DBG_R18_DATA,
				DBG_R19_DATA,
				DBG_R20_DATA,
				DBG_R21_DATA,
				DBG_R22_DATA,
				DBG_R23_DATA,
				DBG_R24_DATA,
				DBG_R25_DATA,
				DBG_R26_DATA,
				DBG_R27_DATA,
				DBG_R28_DATA,
				DBG_R29_DATA,
				DBG_R30_DATA,
				DBG_R31_DATA
	);

	-- Unidade de Controle
	CONTROL0: CONTROL PORT MAP(
				-- in
				CLOCK,
				INSTRUCAO_ID,
				-- out
				RegWrite_ID, 
				ALUSrc_ID,
				ALUOp_ID,
				RegDst_ID,
				MemWrite_ID,
				MemRead_ID,
				MemtoReg_ID,
				Branch_ID,
				OPCODE_ID, 
				FUNCT_ID,
				RD_ADDR_ID,
				RS_ADDR_ID,
				RT_ADDR_ID,
				AddSrc_ID,
				Jump_ID,
				ImmedOrReg_ID
	);
	
	-- REG PIPELINE ID/EX
	RegistradorID_EX0: RegistradorID_EX PORT MAP(
				-- in
				RS_DATA_ID, 
				RT_DATA_ID, 
				IMMED_EXT_ID,
				RD_ADDR_ID,
				PC_ID,
				OPCODE_ID,
				CLOCK,				
				FUNCT_ID,
				-- out
				RS_DATA_EX,
				RT_DATA_EX,
				IMMED_EXT_EX,
				RD_ADDR_EX,
				OPCODE_EX,
				PC_EX,
				FUNCT_EX);
			
	
	-- REG EX ID
	RegistradorEX_0: RegistradorEX PORT MAP(
				-- in
				ALUSrc_ID,
				ALUOp_ID,		
				RegDst_ID,
				CLOCK,
				AddSrc_ID,
				ImmedOrReg_ID,
				-- out
				ALUSrc_EX,	
				ALUOp_EX,	
				RegDST_EX,
				AddSrc_EX,
				ImmedOrReg_EX	
	);
	
	
	-- REG MEM ID
	RegistradorMEM_0: RegistradorMEM PORT MAP(
				-- in
				MemWrite_ID,
				MemRead_ID,
				Branch_ID,
				CLOCK,
				Jump_ID,
				-- out
				MemWrite_EX,
				MemRead_EX,
				Branch_EX,
				Jump_EX
	);
	
	-- REG WB ID
	RegistradorWB_0: RegistradorWB PORT MAP(	  
				-- in
				MemToReg_ID,
				RegWrite_ID,
				CLOCK,
				-- out
				MemToReg_EX,
				RegWrite_EX		
	);
	
	
	-------------------------------------------------------------------------------------------
	-- EX 3
	
	-- MUX ALU SOURCE
	MUXALU0: MUX32_2_1 PORT MAP(
				-- in
				RT_DATA_EX,
				IMMED_EXT_EX,				
				ALUSrc_EX,
				-- out
				ALU_B_EX				
	);	
	
	-- MUX Add SOURCE
	MUXADDER0: MUX32_2_1 PORT MAP(
				-- in
				PC_EX,
				"00000000000000000000000000000000",				
				AddSrc_EX,
				-- out
				ADDER_A_EX				
	);	
		
	-- ADDER (CALC BRANCH)
	ADDERBRANCH0: ADDER PORT MAP(	
				-- in
				ADDER_A_EX, 
				IMMED_EXT_EX,	
				-- out
				SOMADOR_TMP_EX
	);
	
	-- MUX Immed Or Reg
	MUXIMMEDORREG0: MUX32_2_1 PORT MAP(
				-- in
				SOMADOR_TMP_EX,
				RS_DATA_EX,				
				ImmedOrReg_EX,
				-- out
				SOMADOR_EX				
	);	
	
	-- ALU CONTROL	
	ALUControl0: ALUControl PORT MAP(
				-- in
				FUNCT_EX,
				ALUOp_EX,
				OPCODE_EX,
				-- out
				OPERACAO_ALU_EX
	);
	
	ALU0: ALU PORT MAP(
				-- in
				RS_DATA_EX,
				ALU_B_EX,
				OPERACAO_ALU_EX,
				-- out
				ALUResult_EX,
				ZERO_EX
	);
	
	
	-- REG PIPELINE EX/MEM
	RegistradorEX_MEM0: RegistradorEX_MEM PORT MAP(
				-- in
				SOMADOR_EX,
				ZERO_EX,
				ALUResult_EX,
				RT_DATA_EX,
				RD_ADDR_EX,
				CLOCK,
				-- out
				SOMADOR_MEM,
				ZERO_MEM,
				ALUResult_MEM,
				RT_DATA_MEM,
				RD_ADDR_MEM
	);
	
	
	-- REG MEM EX
	RegistradorMEM_1: RegistradorMEM PORT MAP(
				-- in
				MemWrite_EX,
				MemRead_EX,
				Branch_EX,
				CLOCK,
				Jump_EX,
				-- out
				MemWrite_MEM,
				MemRead_MEM,
				Branch_MEM,
				Jump_MEM
	);
	
	-- REG WB EX
	RegistradorWB_1: RegistradorWB PORT MAP(	  
				-- in
				MemToReg_EX,
				RegWrite_EX,
				CLOCK,
				-- out
				MemToReg_MEM,
				RegWrite_MEM		
	);
		
	-------------------------------------------------------------------------------------------
	-- MEM 4

	-- DATA MEMORY
	DATAMEMORY0: DATAMEMORY PORT MAP(	
				-- in
				CLOCK, 
				MemWrite_MEM, 
				MemRead_MEM,
				ALUResult_MEM, 
				RT_DATA_MEM,
				-- out
				MEMREAD_DATA_MEM,
				DBG_MEM0,
				DBG_MEM1,
				DBG_MEM2,
				DBG_MEM3,
				DBG_MEM4,
				DBG_MEM5,
				DBG_MEM6,
				DBG_MEM7
	);	
	
	-- PCSource
	PCSource_MEM <= (Branch_MEM AND ZERO_MEM) OR Jump_MEM;
	
	-- REG PIPELINE MEM/WB
	RegistradorMEM_WB0: RegistradorMEM_WB PORT MAP(
				MEMREAD_DATA_MEM,
				ALUResult_MEM,
				RD_ADDR_MEM,
				CLOCK,
				-- out
				MEMREAD_DATA_WB,
				ALUResult_WB,
				RD_ADDR_WB
	);
	
	-- REG WB MEM
	RegistradorWB_2: RegistradorWB PORT MAP(	 	
				-- in
				MemToReg_MEM,
				RegWrite_MEM,
				CLOCK,				
				-- out
				MemToReg_WB,
				RegWrite_WB		
	);
	
	-------------------------------------------------------------------------------------------
	-- WB	5
	
	-- MemToReg MUX
	MUXMEMTOREG: MUX32_2_1 PORT MAP(
				-- in
				ALUResult_WB,
				MEMREAD_DATA_WB,
				MemToReg_WB,
				-- out
				RegWriteData_WB	
	);	

	-------------------------------------------------------------------------------------------
	-- DBG
	
	DBG_PC_IF <= PC_IF;
	--DBG_PC_ID <= PC_ID;
	DBG_INSTRUCAO_IF <= INSTRUCAO_IF;
	--DBG_INSTRUCAO_ID <= INSTRUCAO_ID;

	--DBG_RegWrite_WB <= RegWrite_WB;
	--DBG_RD_ADDR_WB <= RD_ADDR_WB;
	--DBG_RegWriteData_WB <= RegWriteData_WB;
	--DBG_MEMREAD_DATA_WB <= MEMREAD_DATA_WB;
	--DBG_ALUResult_WB <= ALUResult_WB;
	--DBG_MemToReg_WB <= MemToReg_WB;
			
	
	--DBG_REGWRITE_ID <= RegWrite_ID;
	--DBG_REGWRITE_EX <= RegWrite_EX;
	--DBG_REGWRITE_MEM <= RegWrite_MEM;
	
	--DBG_RS_DATA_ID <= RS_DATA_ID;
	--DBG_RT_DATA_ID <= RT_DATA_ID;
	
	--DBG_RS_DATA_EX <= RS_DATA_EX;
	--DBG_RT_DATA_EX <= RT_DATA_EX;
	
	--DBG_RS_ADDR_ID <= RS_ADDR_ID;
	--DBG_RT_ADDR_ID <= RT_ADDR_ID;
	
	--DBG_OPERACAO_ALU_EX <= OPERACAO_ALU_EX;
	--DBG_FUNCT_EX <= FUNCT_EX;
	
	--DBG_MemWrite_MEM <= MemWrite_MEM; 
	--DBG_MemRead_MEM <= MemRead_MEM;
	--DBG_ALUResult_MEM <= ALUResult_MEM; 
	--DBG_RT_DATA_MEM <= RT_DATA_MEM;
	
	--DBG_Branch_MEM <= Branch_MEM ;
	--DBG_ZERO_MEM <= ZERO_MEM;
	--DBG_SOMADOR_MEM <= SOMADOR_MEM;
	
END ARCHITECTURE ; -- arch